library verilog;
use verilog.vl_types.all;
entity LAB5_121220307_mul_cpu_vlg_tst is
end LAB5_121220307_mul_cpu_vlg_tst;
