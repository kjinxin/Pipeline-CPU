// 指令存储器
module InstructionMemery
(
	input [31:0] addr,   //the address of the IR that we want 
	output [31:0] IR     //  the IR
);
reg [7:0] mem[255:0];

initial begin
	$readmemb("testcode", mem); // 用文件 testcode 初始化 mem
end

/*
initial
begin
	{mem[  3], mem[  2], mem[  1], mem[  0]} <= 32'b001111_00000_01000_00010010_00110100;   // lui	$8, 0x1234
	{mem[  7], mem[  6], mem[  5], mem[  4]} <= 32'b001001_01000_00100_01010000_00000000;   // addiu	$4, $8, 0x5000	#4<=0x12345000
	{mem[ 11], mem[ 10], mem[  9], mem[  8]} <= 32'b001111_00000_01001_01000011_00100001;   // lui	$9, 0x4321
	{mem[ 15], mem[ 14], mem[ 13], mem[ 12]} <= 32'b001000_01001_00101_01010000_00000000;   // addi	$5, $9, 0x5000	#5<=0x43215000
	{mem[ 19], mem[ 18], mem[ 17], mem[ 16]} <= 32'b000000_10000_10000_00110_00000_100000;  // add	$6, $16, $16  # overflow!
	{mem[ 23], mem[ 22], mem[ 21], mem[ 20]} <= 32'b000000_10000_10000_00110_00000_100001;  // addu	$6, $16, $16  # $6=0xEA000000
	{mem[ 27], mem[ 26], mem[ 25], mem[ 24]} <= 32'b000000_00100_00101_00110_00000_100000;  // add	$6, $4, $5  # $6=5555a000
	{mem[ 31], mem[ 30], mem[ 29], mem[ 28]} <= 32'b000000_00100_00101_00110_00000_100010;  // sub	$6, $4, $5  # $6=cf130000
	{mem[ 35], mem[ 34], mem[ 33], mem[ 32]} <= 32'b000000_00100_00101_00110_00000_100011;  // subu	$6, $4, $5  # $6=cf130000
	{mem[ 39], mem[ 38], mem[ 37], mem[ 36]} <= 32'b001000_00000_00111_10101011_11001101;   // addi	$7, $0, 0xabcd
	{mem[ 43], mem[ 42], mem[ 41], mem[ 40]} <= 32'b01111100000001110011110000100000;       // seb 	$7, $7   #ffffffcd
	{mem[ 47], mem[ 46], mem[ 45], mem[ 44]} <= 32'b00111000111001111111000011110000;       // xori	$7, $7, 0xf0f0 ##ffff0f3d
	{mem[ 51], mem[ 50], mem[ 49], mem[ 48]} <= 32'b01110000111000000010000000100001;       // clo	$4, $7  # $4 = 16
	{mem[ 55], mem[ 54], mem[ 53], mem[ 52]} <= 32'b01110000100000000011100000100000;       // clz	$7, $4  # $7 = 27
	{mem[ 59], mem[ 58], mem[ 57], mem[ 56]} <= 32'b000000_00000_10001_01010_10000_000011;  // sra $10, $17, 16 ## $10=$17 >>a 16
	{mem[ 63], mem[ 62], mem[ 61], mem[ 60]} <= 32'b000000_00100_10001_01010_00000_000111;  // srav $10, $17, $4 ## $10=$17 >>a 16
	{mem[ 67], mem[ 66], mem[ 65], mem[ 64]} <= 32'b000000_00000_10001_01010_10000_000000;  // sll $10, $17, 16 ## $10=$17 <<l 16
	{mem[ 71], mem[ 70], mem[ 69], mem[ 68]} <= 32'b000000_00100_10001_01010_00000_000100;  // sllv $10, $17, $4 ## $10=$17 <<l 16
	{mem[ 75], mem[ 74], mem[ 73], mem[ 72]} <= 32'b000000_00000_10001_01010_10000_000010;  // srl $10, $17, 16 ## $10=$17 >>l 16
	{mem[ 79], mem[ 78], mem[ 77], mem[ 76]} <= 32'b000000_00100_10001_01010_00000_000110;  // srlv $10, $17, $4 ## $10=$17 >>l 16
	{mem[ 83], mem[ 82], mem[ 81], mem[ 80]} <= 32'b000000_00001_00101_00101_00100_000010;  // rotr	$5, $5, 4    # $5=0x04321500
	{mem[ 87], mem[ 86], mem[ 85], mem[ 84]} <= 32'b000000_00100_00101_00101_00001_000110;  // rotrv  $5, $5, $4   # $5=0x15000432
	{mem[ 91], mem[ 90], mem[ 89], mem[ 88]} <= 32'b00100101000001000101011001111000;       // addiu	$4, $8, 0x5678	# $4<=0x12345678
	{mem[ 95], mem[ 94], mem[ 93], mem[ 92]} <= 32'b000000_00100_00101_00110_00000_100111;  // nor	$6, $4, $5
	{mem[ 99], mem[ 98], mem[ 97], mem[ 96]} <= 32'b000000_00100_00101_00110_00000_100100;  // and	$6, $4, $5
	{mem[103], mem[102], mem[101], mem[100]} <= 32'b000000_00100_00101_00110_00000_100101;  // or 	$6, $4, $5
	{mem[107], mem[106], mem[105], mem[104]} <= 32'b000000_00100_00101_00110_00000_100110;  // xor 	$6, $4, $5
	{mem[111], mem[110], mem[109], mem[108]} <= 32'b001100_00000_00111_10101011_11001101;   // andi	$7, $0, 0xabcd
	{mem[115], mem[114], mem[113], mem[112]} <= 32'b001101_00000_00111_10101011_11001101;   // ori	$7, $0, 0xabcd
	{mem[119], mem[118], mem[117], mem[116]} <= 32'b00111100000010011000001100100001;       // lui	$9, 0x8321
	{mem[123], mem[122], mem[121], mem[120]} <= 32'b00100001001001010101000000000000;       // addi	$5, $9, 0x5000	# $5<=0x83215000
   {mem[127], mem[126], mem[125], mem[124]} <= 32'b00000100101100010000000000001010;       // bgezal $5, +10 # false
	{mem[131], mem[130], mem[129], mem[128]} <= 32'b000000_00100_00101_00110_00000_101010;  // slt  $6, $4, $5  # $6<=0x0
	{mem[135], mem[134], mem[133], mem[132]} <= 32'b000000_00100_00101_00110_00000_101011;  // sltu $6, $4, $5  # $6<=0x1
	{mem[139], mem[138], mem[137], mem[136]} <= 32'b00000000101001000011000000101011;       // sltu 	$6, $5, $4  # $6<=0x0
	{mem[143], mem[142], mem[141], mem[140]} <= 32'b00101000110001010000000000000010;       // slti	$5, $6, 2 # $5<=0x1
	{mem[147], mem[146], mem[145], mem[144]} <= 32'b00000100101100010000000000000011;       // bgezal $5, +3
	{mem[151], mem[150], mem[149], mem[148]} <= 32'b00000000000000000000000000000000;	     // nop
	{mem[155], mem[154], mem[153], mem[152]} <= 32'b00000000000000000000000000000000;	     // nop
	{mem[159], mem[158], mem[157], mem[156]} <= 32'b00000000000000000000000000000000;	     // nop
	{mem[163], mem[162], mem[161], mem[160]} <= 32'b10101100000001000000000000000000;       // sw  $4, 0($0)
	{mem[167], mem[166], mem[165], mem[164]} <= 32'b10001100000000010000000000000000;       // lw  $1, 0($0)
	{mem[171], mem[170], mem[169], mem[168]} <= 32'b10111000000100010000000000000101;       // swr $17, 5($0) # $17==0xABCD4321
	{mem[175], mem[174], mem[173], mem[172]} <= 32'b10001000000000100000000000000010;       // lwl $2, 2($0)
	{mem[179], mem[178], mem[177], mem[176]} <= 32'b10011000000000100000000000000101;       // lwr $2, 5($0)
	{mem[183], mem[182], mem[181], mem[180]} <= 32'b00000000010000000100100000100000;       // add $9, $2, $0 # $9=$2=0x56784321
	{mem[187], mem[186], mem[185], mem[184]} <= 32'b10101000000100010000000000000010;       // swl $17, 2($0)
	{mem[191], mem[190], mem[189], mem[188]} <= 32'b10001100000000010000000000000000;       // lw  $1, 0($0) # 0x1234ABCD
	{mem[195], mem[194], mem[193], mem[192]} <= 32'b101000_00000_00001_00000000_00000111;   // sb $1, 7($0)  # store byte "CD"
	{mem[199], mem[198], mem[197], mem[196]} <= 32'b100000_00000_00010_00000000_00000111;   // lb $2, 7($0)  # $2 = FFFFFFCD
	{mem[203], mem[202], mem[201], mem[200]} <= 32'b100100_00000_00010_00000000_00000111;   // lbu $2, 7($0) # $2 = 000000CD
	{mem[207], mem[206], mem[205], mem[204]} <= 32'b000000_00001_00000_01001_00000_100000;  // addu $9, $1, $0  # $9=$1=0x1234ABCD
	{mem[211], mem[210], mem[209], mem[208]} <= 32'b101001_00000_00001_00000000_00000111;   // sh $1, 7($0)  # store halfword "ABCD"
	{mem[215], mem[214], mem[213], mem[212]} <= 32'b100001_00000_00010_00000000_00000111;   // lh $2, 7($0)  # $2 = FFFFABCD
	{mem[219], mem[218], mem[217], mem[216]} <= 32'b100101_00000_00010_00000000_00000111;   // lhu $2, 7($0) # $2 = 0000ABCD
	{mem[223], mem[222], mem[221], mem[220]} <= 32'b0;
	{mem[227], mem[226], mem[225], mem[224]} <= 32'b0;
	{mem[231], mem[230], mem[229], mem[228]} <= 32'b0;
	{mem[235], mem[234], mem[233], mem[232]} <= 32'b0;
	{mem[239], mem[238], mem[237], mem[236]} <= 32'b0;
	{mem[243], mem[242], mem[241], mem[240]} <= 32'b0;
	{mem[247], mem[246], mem[245], mem[244]} <= 32'b0;
	{mem[251], mem[250], mem[249], mem[248]} <= 32'b0;
	{mem[255], mem[254], mem[253], mem[252]} <= 32'b000010_000000_000000_000000_000000_00;  // j 0
end
*/
assign IR={mem[addr+3],mem[addr+2],mem[addr+1],mem[addr]};
endmodule 
