library verilog;
use verilog.vl_types.all;
entity lab2_121220307_ARM32_vlg_tst is
end lab2_121220307_ARM32_vlg_tst;
