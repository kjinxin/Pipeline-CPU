library verilog;
use verilog.vl_types.all;
entity lab3_121220307_ARM32_vlg_tst is
end lab3_121220307_ARM32_vlg_tst;
