library verilog;
use verilog.vl_types.all;
entity single_cpu_vlg_tst is
end single_cpu_vlg_tst;
