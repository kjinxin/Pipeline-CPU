library verilog;
use verilog.vl_types.all;
entity lab1_121220307_MIPS4_vlg_tst is
end lab1_121220307_MIPS4_vlg_tst;
